```vhdl
entity counter is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           count : out  UNSIGNED(3 downto 0)); --Corrected to use unsigned type
end entity;

architecture behavioral of counter is
    signal internal_count : UNSIGNED(3 downto 0) := (others => '0');
begin
    process (clk, rst)
    begin
        if rst = '1' then
            internal_count <= (others => '0');
        elsif rising_edge(clk) then
            internal_count <= internal_count + 1;
        end if;
    end process;
    count <= internal_count;
end architecture;
```